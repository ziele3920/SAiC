** Profile: "SCHEMATIC1-symulacja"  [ f:\air\saic\saic\sim-02\rozniczkujacy-schematic1-symulacja.sim ] 

** Creating circuit file "rozniczkujacy-schematic1-symulacja.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 3000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rozniczkujacy-SCHEMATIC1.net" 


.END
