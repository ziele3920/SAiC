** Profile: "SCHEMATIC1-symulacja-filtr"  [ F:\AiR\SAiC\sprawka\SAiC\sim\filtr_sr-SCHEMATIC1-symulacja-filtr.sim ] 

** Creating circuit file "filtr_sr-SCHEMATIC1-symulacja-filtr.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 10 100000
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\filtr_sr-SCHEMATIC1.net" 


.END
