** Profile: "SCHEMATIC1-sp"  [ f:\air\saic\sim\zas-schematic1-sp.sim ] 

** Creating circuit file "zas-schematic1-sp.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\zas-SCHEMATIC1.net" 


.END
