** Profile: "SCHEMATIC1-wzmacniacz2sim"  [ c:\users\jakub\desktop\saic\wzmacniacz2\wzmacniacz2-schematic1-wzmacniacz2sim.sim ] 

** Creating circuit file "wzmacniacz2-schematic1-wzmacniacz2sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 10Meg
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\wzmacniacz2-SCHEMATIC1.net" 


.END
