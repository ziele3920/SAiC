** Profile: "SCHEMATIC1-symulacja-filtr"  [ c:\users\jakub\desktop\saic\saic\sim\filtr_sr-schematic1-symulacja-filtr.sim ] 

** Creating circuit file "filtr_sr-schematic1-symulacja-filtr.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 50 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\filtr_sr-SCHEMATIC1.net" 


.END
