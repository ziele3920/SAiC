** Profile: "SCHEMATIC1-symulacja"  [ F:\AIR\SAiC\projekty\02\rozniczkujacy-SCHEMATIC1-symulacja.sim ] 

** Creating circuit file "rozniczkujacy-SCHEMATIC1-symulacja.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rozniczkujacy-SCHEMATIC1.net" 


.END
